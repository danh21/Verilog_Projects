`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:54:01 12/09/2021 
// Design Name: 
// Module Name:    button 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module button
	#(parameter A = 500000)	//m_tick
	(
	input reset, clk, btn,
	output reg db
    );
	localparam [2:0] 
		zero = 3'b000, wait1_1 = 3'b001, wait1_2 = 3'b010, wait1_3 = 3'b011,
		one = 3'b100, wait0_1 = 3'b101, wait0_2 = 3'b110, wait0_3 = 3'b111;
	localparam N = 19;
// signal declaration
	reg [N-1:0] q_reg;
	wire [N-1:0] q_next;
	wire m_tick;
	reg [2:0] state_reg, state_next;
// counter to generate 10ms tick
always @(posedge clk, posedge reset)
	if (reset)
		q_reg <= 0;
	else
		q_reg <= q_next;
// next state logic
assign q_next = (q_reg == A) ? 0 : q_reg + 1;
// output tick
assign m_tick = (q_reg == 0) ? 1'b1 : 1'b0;
// debouncing FSM
// state register 
always @ (posedge clk, posedge reset)
	if (reset)
		state_reg <= zero;
	else 
		state_reg <= state_next;
// next state logic and output logic
always @*
begin
	state_next = state_reg; // default state
	db = 1'b0;
	case (state_reg)
		zero: if (btn) state_next = wait1_1;
		wait1_1: if (~btn) state_next = zero;
					else 
						if (m_tick) state_next = wait1_2;
		wait1_2: if (~btn) state_next = zero;
					else
						if (m_tick) state_next = wait1_3;
		wait1_3: if (~btn) state_next = zero;
					else
						if (m_tick) state_next = one;
		one: 
		begin
			db = 1'b1;
			if (~btn) state_next = wait0_1;
		end
		wait0_1: 
		begin
			db = 1'b1;
			if (btn)
				state_next = one;
			else
				if (m_tick) state_next = wait0_2;
		end
		wait0_2: 
		begin
			db = 1'b1;
			if (btn)
				state_next = one;
			else
				if (m_tick) state_next = wait0_3;
		end
		wait0_3: 
		begin
			db = 1'b1;
			if (btn)
				state_next = one;
			else
				if (m_tick) state_next = zero;		
		end
		default: state_next = zero;
	endcase
end
endmodule
